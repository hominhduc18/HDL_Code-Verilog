module IC82c19(s,i,e,y);
input [3:0]s;
input i;
input [15:0]e;
output y;
reg y;
always @(*)
begin
if(i==1'b1)
y=1;
else
	begin 
		case(s)
		4'b0000:y=~e[0];
		4'b0001:y=~e[1];
		4'b0010:y=~e[2];
		4'b0011:y=~e[3];
		4'b0100:y=~e[4];
      4'b0101:y=~e[5];
		4'b0110:y=~e[6];
		4'b0111:y=~e[7];
		4'b1000:y=~e[8];
		4'b1001:y=~e[9];
		4'b1010:y=~e[10];
		4'b1011:y=~e[11];
		4'b1100:y=~e[12];
		4'b1101:y=~e[13];
		4'b1110:y=~e[14];
		4'b1111:y=~e[15];
		endcase
	end
end 
endmodule

module TB_IC82c19();
reg [3:0]s;
reg [15:0]e;
reg i;
wire y;
initial 
begin 
i=0;
s=4'b0000;
e=16'b0000000000000001;
#100
i=0;
s=4'b0001;
e=16'b0000000000000010;
#100
i=0;
s=4'b0010;
e=16'b0000000000000100;
#100
i=0;
s=4'b0011;
e=16'b0000000000001000;
#100
i=0;
s=4'b0100;
e=16'b0000000000010000;
#100
i=0;
s=4'b0101;
e=16'b0000000000100000;
#100
i=0;
s=4'b0110;
e=16'b0000000001000000;
#100
i=0;
s=4'b0111;
e=16'b0000000010000000;
#100
i=0;
s=4'b1000;
e=16'b0000000100000000;
#100
i=0;
s=4'b1001;
e=16'b0000001000000000;
#100
i=0;
s=4'b1010;
e=16'b0000010000000000;
#100
i=0;
s=4'b1011;
e=16'b0000100000000000;
#100
i=0;
s=4'b1100;
e=16'b0001000000000000;
#100
i=0;
s=4'b1101;
e=16'b0010000000000000;
#100
i=0;
s=4'b1110;
e=16'b0100000000000000;
#100
i=0;
s=4'b1111;
e=16'b1000000000000000;
#100
i=0;
s=4'b0000;
e=16'b111111111111110;
#100
i=0;
s=4'b0001;
e=16'b1111111111111101;
#100
i=0;
s=4'b0010;
e=16'b1111111111111011;
#100
i=0;
s=4'b0011;
e=16'b1111111111110111;
#100
i=0;
s=4'b0100;
e=16'b1111111111101111;
#100
i=0;
s=4'b0101;
e=16'b1111111111011111;
#100
i=0;
s=4'b0110;
e=16'b1111111110111111;
#100
i=0;
s=4'b0111;
e=16'b1111111101111111;
#100
i=0;
s=4'b1000;
e=16'b1111111011111111;
#100
i=0;
s=4'b1001;
e=16'b1111110111111111;
#100
i=0;
s=4'b1010;
e=16'b1111101111111111;
#100
i=0;
s=4'b1011;
e=16'b1111011111111111;
#100
i=0;
s=4'b1100;
e=16'b1110111111111111;
#100
i=0;
s=4'b1101;
e=16'b1101111111111111;
#100
i=0;
s=4'b1110;
e=16'b1011111111111111;
#100
i=0;
s=4'b1111;
e=16'b0111111111111111;
#3500 $finish;
end
IC82c19 D(.s(s),.i(i),.e(e),.y(y));
endmodule
