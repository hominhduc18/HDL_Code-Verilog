module bai10(A,Y);
input [4:0]A;
output Y;
reg Y;
always @(*)
begin 
if((A%2!=0 && A>=2 && A%3!=0) || (A==2 || A==3))
Y=1'b1;
else
Y=1'b0;
end
endmodule
module TB_bai10();
reg [4:0]A;
wire Y;
initial
begin
A = 5'b00000; 
#100
A = 5'b00001;
#100
A = 5'b00010; 
#100
A = 5'b00011;
#100
A = 5'b00100;
#100
A = 5'b00101;
#100
A = 5'b00110;
#100
A=5'b00111;
#100
A = 5'b01000;
#100
A = 5'b01001; 
#100
A = 5'b01010;
#100
A = 5'b01011;
#100
A = 5'b01100;
#100
A = 5'b01101;
#100
A = 5'b01110;
#100
A = 5'b01111; 
#100
A = 5'b10000;
#100
A = 5'b10001;
#100
A = 5'b10010;
#100
A = 5'b10011;
#100
A=5'b10100;
#100
A = 5'b10101;
#100
A = 5'b10110; 
#100
A = 5'b10111;
#100
A = 5'b11000;
#100
A = 5'b11001;
#100
A = 5'b11010;
#100
A=5'b11011;
#100
A = 5'b11100;
#100
A = 5'b11101; 
#100
A = 5'b11110;
#100
A = 5'b11111;
#5000 $finish;
end
bai10 D(.A(A),.Y(Y));
endmodule

